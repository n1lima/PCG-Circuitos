module xor (a, b, s);
    input a;       
    input b;       
    output y;       

    assign s = a ^ b;

endmodule
